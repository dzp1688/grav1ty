`default_nettype none

package obu_parser_pkg;
    localparam PARSER_DATA_WIDTH = 32;
endpackage

