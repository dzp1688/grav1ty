`default_nettype none

package obu_parser_pkg;
    localparam PARSER_DATA_WIDTH = 32;
    localparam PAD_LEN_WIDTH = $clog2(PARSER_DATA_WIDTH) + 1;
endpackage

