`default_nettype none

module field_aligner ()

endmodule
